//sample module

module buffer(input a,output reg y);

always@(a)
y=a;

endmodule